

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 256;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr[30:2] < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin

			ROMDATA[0] <= 32'b00001000000000000000000000000100;	//RESET:	j	INIT
			ROMDATA[1] <= 32'b00001000000000000000000001100011;	//ILLOP:	j	INTRPT
			ROMDATA[2] <= 32'b00001000000000000000000000000011;	//XADR:	j	EXPT
			ROMDATA[3] <= 32'b00000011111000000000000000001000;	//EXPT:	jr	$ra
			ROMDATA[4] <= 32'b00100000000010000000000000111111;	//INIT:	addi	$t0,	$zero,	0x3f	#0
			ROMDATA[5] <= 32'b10101100000010000000000000000000;	//	sw	$t0,	0($zero)
			ROMDATA[6] <= 32'b00100000000010010000000000000110;	//	addi	$t1,	$zero,	0x06	#1
			ROMDATA[7] <= 32'b10101100000010010000000000000100;	//	sw	$t1,	4($zero)
			ROMDATA[8] <= 32'b00100000000010000000000001011011;	//	addi	$t0,	$zero,	0x5b	#2
			ROMDATA[9] <= 32'b10101100000010000000000000001000;	//	sw	$t0,	8($zero)
			ROMDATA[10] <= 32'b00100000000010010000000001001111;	//	addi	$t1,	$zero,	0x4f	#3
			ROMDATA[11] <= 32'b10101100000010010000000000001100;	//	sw	$t1,	12($zero)
			ROMDATA[12] <= 32'b00100000000010000000000001100110;	//	addi	$t0,	$zero,	0x66	#4
			ROMDATA[13] <= 32'b10101100000010000000000000010000;	//	sw	$t0,	16($zero)
			ROMDATA[14] <= 32'b00100000000010010000000001101101;	//	addi	$t1,	$zero,	0x6d	#5
			ROMDATA[15] <= 32'b10101100000010010000000000010100;	//	sw	$t1,	20($zero)
			ROMDATA[16] <= 32'b00100000000010000000000001111101;	//	addi	$t0,	$zero,	0x7d	#6
			ROMDATA[17] <= 32'b10101100000010000000000000011000;	//	sw	$t0,	24($zero)
			ROMDATA[18] <= 32'b00100000000010010000000000000111;	//	addi	$t1,	$zero,	0x07	#7
			ROMDATA[19] <= 32'b10101100000010010000000000011100;	//	sw	$t1,	28($zero)
			ROMDATA[20] <= 32'b00100000000010000000000001111111;	//	addi	$t0,	$zero,	0x7f	#8
			ROMDATA[21] <= 32'b10101100000010000000000000100000;	//	sw	$t0,	32($zero)
			ROMDATA[22] <= 32'b00100000000010010000000001101111;	//	addi	$t1,	$zero,	0x6f	#9
			ROMDATA[23] <= 32'b10101100000010010000000000100100;	//	sw	$t1,	36($zero)
			ROMDATA[24] <= 32'b00100000000010000000000001110111;	//	addi	$t0,	$zero,	0x77	#a
			ROMDATA[25] <= 32'b10101100000010000000000000101000;	//	sw	$t0,	40($zero)
			ROMDATA[26] <= 32'b00100000000010010000000001111100;	//	addi	$t1,	$zero,	0x7c	#b
			ROMDATA[27] <= 32'b10101100000010010000000000101100;	//	sw	$t1,	44($zero)
			ROMDATA[28] <= 32'b00100000000010000000000000111001;	//	addi	$t0,	$zero,	0x39	#c
			ROMDATA[29] <= 32'b10101100000010000000000000110000;	//	sw	$t0,	48($zero)
			ROMDATA[30] <= 32'b00100000000010010000000001011110;	//	addi	$t1,	$zero,	0x5e	#d
			ROMDATA[31] <= 32'b10101100000010010000000000110100;	//	sw	$t1,	52($zero)
			ROMDATA[32] <= 32'b00100000000010000000000001111011;	//	addi	$t0,	$zero,	0x7b	#e
			ROMDATA[33] <= 32'b10101100000010000000000000111000;	//	sw	$t0,	56($zero)
			ROMDATA[34] <= 32'b00100000000010010000000001110001;	//	addi	$t1,	$zero,	0x71	#f
			ROMDATA[35] <= 32'b10101100000010010000000000111100;	//	sw	$t1,	60($zero)
			ROMDATA[36] <= 32'b00100000000101110000000000000001;	//	addi	$s7,	$zero,	1	#digi
			ROMDATA[37] <= 32'b00111100000111000100000000000000;	//	lui	$gp,	0x4000
			ROMDATA[38] <= 32'b10101111100000000000000000001000;	//	sw	$zero,	8($gp)		#set Timer COntrol
			ROMDATA[39] <= 32'b00100000000010010000000000000011;	//	addi	$t1,	$zero,	3
			ROMDATA[40] <= 32'b10101111100010010000000000100000;	//	sw	$t1,	32($gp)		#set UART Control
			ROMDATA[41] <= 32'b00001000000000000000000000101001;	//STAY:	j	STAY			#stay here in the end
			ROMDATA[42] <= 32'b00111100000011011111111111111111;	//MAIN:	lui	$t5,	0xffff
			ROMDATA[43] <= 32'b00110101101011010011110010101111;	//	ori	$t5,	0x3caf
			ROMDATA[44] <= 32'b10101111100011010000000000000000;	//	sw	$t5,	0($gp)
			ROMDATA[45] <= 32'b10101111100011010000000000000100;	//	sw	$t5,	4($gp)
			ROMDATA[46] <= 32'b00100000000011100000000000000011;	//	addi	$t6,	$zero,	3
			ROMDATA[47] <= 32'b10101111100011100000000000001000;	//	sw	$t6,	8($gp)
			ROMDATA[48] <= 32'b00100011101111011111111111110000;	//bgcd:	addi	$sp,	$sp,	-16
			ROMDATA[49] <= 32'b10101111101101000000000000001100;	//	sw	$s4,	12($sp)		#counter of 2
			ROMDATA[50] <= 32'b10101111101100100000000000001000;	//	sw	$s2,	8($sp)		#num1even
			ROMDATA[51] <= 32'b10101111101100110000000000000100;	//	sw	$s3,	4($sp)		#num2even
			ROMDATA[52] <= 32'b10101111101111110000000000000000;	//	sw	$ra,	0($sp)
			ROMDATA[53] <= 32'b00010000100000000000000000100001;	//	beq	$a0,	$zero,	Return1	#num1==0
			ROMDATA[54] <= 32'b00010000101000000000000000100010;	//	beq	$a1,	$zero,	Return2	#num2==0
			ROMDATA[55] <= 32'b00100000000010010000000000000001;	//	addi	$t1,	$zero,	1
			ROMDATA[56] <= 32'b00000000100010011001000000100100;	//	and	$s2,	$a0,	$t1	#num1even
			ROMDATA[57] <= 32'b00000000101010011001100000100100;	//	and	$s3,	$a1,	$t1	#num2even
			ROMDATA[58] <= 32'b00100000000010010000000000000001;	//	addi	$t1,	$zero,	1
			ROMDATA[59] <= 32'b00000010010100110101000000100101;	//	or	$t2,	$s2,	$s3
			ROMDATA[60] <= 32'b00010101001010100000000000000100;	//	bne	$t1,	$t2,	ALLEVEN
			ROMDATA[61] <= 32'b00000010010100110100100000100100;	//	and	$t1,	$s2,	$s3
			ROMDATA[62] <= 32'b00010101001000000000000000001100;	//	bne	$t1,	$zero,	ALLODD
			ROMDATA[63] <= 32'b00010010010000000000000000000101;	//	beq	$s2,	$zero,	ONEEVEN
			ROMDATA[64] <= 32'b00010010011000000000000000000111;	//	beq	$s3,	$zero,	TWOEVEN
			ROMDATA[65] <= 32'b00000000000001000010000001000010;	//ALLEVEN:srl	$a0,	$a0,	1	# num1 = num1 >> 1
			ROMDATA[66] <= 32'b00000000000001010010100001000010;	//    	srl	$a1,	$a1,	1	# num2 = num2 >> 1
			ROMDATA[67] <= 32'b00100010100101000000000000000001;	//    	addi	$s4,	$s4,	1	# s4++
			ROMDATA[68] <= 32'b00001100000000000000000000110000;	//    	jal	bgcd
			ROMDATA[69] <= 32'b00000000000001000010000001000010;	//ONEEVEN:srl	$a0,	$a0,	1		#num1 = num1>>1
			ROMDATA[70] <= 32'b00000000101000000010100000100000;	//	add	$a1,	$a1,	$zero	#num2 keep
			ROMDATA[71] <= 32'b00001100000000000000000000110000;	//	jal	bgcd
			ROMDATA[72] <= 32'b00000000000001010010100001000010;	//TWOEVEN:srl	$a1,	$a1,	1		#num2 = num2>>1
			ROMDATA[73] <= 32'b00000000100000000010000000100000;	//	add	$a0,	$a0,	$zero	#num1 keep
			ROMDATA[74] <= 32'b00001100000000000000000000110000;	//	jal 	bgcd
			ROMDATA[75] <= 32'b00000000100001010100100000101010;	//ALLODD:	slt	$t1,	$a0,	$a1	#num1<num2 -> t1=1
			ROMDATA[76] <= 32'b00010101001000000000000000000101;	//	bne	$t1,	$zero,	ONELTWO
			ROMDATA[77] <= 32'b00000000100001010100100000100010;	//	sub	$t1,	$a0,	$a1	#num1>num2
			ROMDATA[78] <= 32'b00000000000010010100100001000010;	//	srl	$t1,	$t1,	1
			ROMDATA[79] <= 32'b00000001001000000010000000100000;	//	add	$a0	$t1,	$zero	#num1 = (num1 - num2)>>1
			ROMDATA[80] <= 32'b00000000101000000010100000100000;	//	add	$a1,	$a1,	$zero	#num2 keep
			ROMDATA[81] <= 32'b00001100000000000000000000110000;	//	jal	bgcd
			ROMDATA[82] <= 32'b00000000101001000100100000100010;	//ONELTWO:sub	$t1,	$a1,	$a0	#num1<num2
			ROMDATA[83] <= 32'b00000000000010010100100001000010;	//	srl	$t1,	$t1,	1
			ROMDATA[84] <= 32'b00000001001000000010100000100000;	//	add	$a1,	$t1,	$zero	#num2 = (num2 - num1)>>1;
			ROMDATA[85] <= 32'b00000000100000000010000000100000;	//	add	$a0,	$a0,	$zero	#num1 keep
			ROMDATA[86] <= 32'b00001100000000000000000000110000;	//	jal	bgcd
			ROMDATA[87] <= 32'b00000000000001010001000000100000;	//Return1:add	$v0,	$zero,	$a1	#num1==0 #return num2
			ROMDATA[88] <= 32'b00001000000000000000000001011011;	//	j	LOOP
			ROMDATA[89] <= 32'b00000000000001000001000000100000;	//Return2:add	$v0,	$zero,	$a0	#num2==0 #return num1
			ROMDATA[90] <= 32'b00001000000000000000000001011011;	//	j	LOOP
			ROMDATA[91] <= 32'b00010010100000000000000000000100;	//LOOP:	beq	$s4,	$zero,	GCDFIN
			ROMDATA[92] <= 32'b00000000000000100001000001000000;	//	sll	$v0,	$v0,	1
			ROMDATA[93] <= 32'b00100000000010010000000000000001;	//	addi	$t1,	$zero,	1
			ROMDATA[94] <= 32'b00000010100010011010000000100010;	//	sub	$s4,	$s4,	$t1
			ROMDATA[95] <= 32'b00001000000000000000000001011011;	//	j	LOOP
			ROMDATA[96] <= 32'b10101111100000100000000000011000;	//GCDFIN:	sw	$v0,	24($gp)
			ROMDATA[97] <= 32'b10101111100000100000000000001100;	//	sw	$v0,	12($gp)
			ROMDATA[98] <= 32'b00001000000000000000000000101001;	//	j	STAY
			ROMDATA[99] <= 32'b10001111100011110000000000100000;	//INTRPT:	lw	$t7,	32($gp)		#Load UART Control
			ROMDATA[100] <= 32'b00101001111010010000000000001000;	//	slti	$t1,	$t7,	8	#Judge whether is sending intrpt
			ROMDATA[101] <= 32'b00010101001000000000000000001110;	//	bne	$t1,	$zero,	TIMER
			ROMDATA[102] <= 32'b10001111100100000000000000011100;	//	lw	$s0,	28($gp)
			ROMDATA[103] <= 32'b00010110110000000000000000000100;	//	bne	$s6,	$zero,	ALREADY	#Judge whether has already gotten a parameter
			ROMDATA[104] <= 32'b00000000000100000010000000100000;	//	add	$a0,	$zero,	$s0
			ROMDATA[105] <= 32'b00000000000100001100000000100000;	//	add $t8,	$zero,	$s0
			ROMDATA[106] <= 32'b00100010110101100000000000000001;	//	addi	$s6,	$s6,	1
			ROMDATA[107] <= 32'b00000011010000000000000000001000;	//	jr	$k0
			ROMDATA[108] <= 32'b00000000000100000010100000100000;	//ALREADY:add	$a1,	$zero,	$s0
			ROMDATA[109] <= 32'b00000000000100001100100000100000;	//	add	$t9,	$zero,	$s0
			ROMDATA[110] <= 32'b00000000000000001011000000100000;	//	add	$s6,	$zero,	$zero
			ROMDATA[111] <= 32'b00000000000000001000000000100000;	//	add	$s0,	$zero,	$zero
			ROMDATA[112] <= 32'b00100000000010010000000000000001;	//	addi	$t1,	$zero,	1
			ROMDATA[113] <= 32'b10101111100010010000000000100000;	//	sw	$t1,	32($gp)
			ROMDATA[114] <= 32'b00100011010110100000000000000100;	//	addi	$k0,	$k0,	4
			ROMDATA[115] <= 32'b00000011010000000000000000001000;	//	jr	$k0
			ROMDATA[116] <= 32'b00111100000010001111111111111111;	//TIMER:	lui	$t0,	0xffff
			ROMDATA[117] <= 32'b00110101000010001111111111111001;	//	ori	$t0,	$t0,	0xfff9
			ROMDATA[118] <= 32'b10001111100010010000000000001000;	//	lw	$t1,	8($gp)
			ROMDATA[119] <= 32'b00000001001010000100100000100100;	//	and	$t1,	$t1,	$t0
			ROMDATA[120] <= 32'b10101111100010010000000000001000;	//	sw	$t1,	8($gp)
			ROMDATA[121] <= 32'b00000000000101110101001000000000;	//DIGI:	sll	$t2,	$s7,	8
			ROMDATA[122] <= 32'b00101001010011110000010000000000;	//	slti	$t7,	$t2,	0x400
			ROMDATA[123] <= 32'b00010101111000000000000000000111;	//	bne	$t7,	$zero,	SECOND
			ROMDATA[124] <= 32'b00101001010011100000100000000000;	//FIRST:	slti	$t6,	$t2,	0x800
			ROMDATA[125] <= 32'b00010101110000000000000000000011;	//	bne	$t6,	$zero	FIRSTL
			ROMDATA[126] <= 32'b00110011000011000000000011110000;	//FIRSTH:	andi	$t4,	$t8,	0x00f0
			ROMDATA[127] <= 32'b00000000000011000110000100000010;	//	srl	$t4,	$t4,	4
			ROMDATA[128] <= 32'b00001000000000000000000010001001;	//	j	DISPLAY
			ROMDATA[129] <= 32'b00110011000011000000000000001111;	//FIRSTL:	andi	$t4,	$t8,	0x000f
			ROMDATA[130] <= 32'b00001000000000000000000010001001;	//	j	DISPLAY
			ROMDATA[131] <= 32'b00101001010011100000001000000000;	//SECOND:	slti 	$t6,	$t2,	0x200
			ROMDATA[132] <= 32'b00010101110000000000000000000011;	//	bne	$t6,	$zero,	SECONDL
			ROMDATA[133] <= 32'b00110011001011000000000011110000;	//SECONDH:andi	$t4,	$t9,	0x00f0
			ROMDATA[134] <= 32'b00000000000011000110000100000010;	//	srl	$t4,	$t4,	4
			ROMDATA[135] <= 32'b00001000000000000000000010001001;	//	j	DISPLAY
			ROMDATA[136] <= 32'b00110011001011000000000000001111;	//SECONDL:andi	$t4,	$t9,	0x000f
			ROMDATA[137] <= 32'b00000000000011000110000010000000;	//DISPLAY:sll	$t4,	$t4,	2
			ROMDATA[138] <= 32'b10001101100011000000000000000000;	//	lw	$t4,	0($t4)
			ROMDATA[139] <= 32'b00000001010011000101000000100000;	//	add	$t2,	$t2,	$t4
			ROMDATA[140] <= 32'b10101111100010100000000000010100;	//	sw	$t2,	20($gp)
			ROMDATA[141] <= 32'b00000000000101111011100001000000;	//	sll	$s7,	$s7,	1
			ROMDATA[142] <= 32'b00101010111011100000000000001001;	//	slti	$t6,	$s7,	0x09
			ROMDATA[143] <= 32'b00010101110000000000000000000001;	//	bne	$t6,	$zero,	FIN
			ROMDATA[144] <= 32'b00100000000101110000000000000001;	//	addi	$s7,	$zero,	1
			ROMDATA[145] <= 32'b10001111100010010000000000001000;	//FIN:	lw	$t1,	8($gp)
			ROMDATA[146] <= 32'b00110101001010010000000000000010;	//	ori	$t1,	$t1,	0x0002
			ROMDATA[147] <= 32'b10101111100010010000000000001000;	//	sw	$t1,	8($gp)
			ROMDATA[148] <= 32'b00000011010000000000000000001000;	//	jr	$k0


		for (i=149;i<ROM_SIZE;i=i+1) begin
			ROMDATA[i] <= 32'b0;
		end
end
endmodule
